------------------------------------------
-----------COMANDOS PARA LCD--------------
------------�NO MODIFICAR!---------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;

package COMANDOS_LCDSPI_REVA is

FUNCTION LCD_INI(DATO : STD_LOGIC_VECTOR(1 DOWNTO 0)) RETURN STD_LOGIC_VECTOR;
FUNCTION CHAR(DATO1 : INTEGER) RETURN STD_LOGIC_VECTOR;
FUNCTION POS(DATO2,DATO3 : INTEGER) RETURN STD_LOGIC_VECTOR;
FUNCTION CHAR_ASCII(DATO6 : STD_LOGIC_VECTOR(7 DOWNTO 0))RETURN STD_LOGIC_VECTOR;
FUNCTION CODIGO_FIN(DATO7 : INTEGER) RETURN STD_LOGIC_VECTOR;
FUNCTION BUCLE_INI(DATO8 : INTEGER)RETURN STD_LOGIC_VECTOR;
FUNCTION BUCLE_FIN(DATO9 : INTEGER)RETURN STD_LOGIC_VECTOR;
FUNCTION INT_NUM(DATO10 : INTEGER)RETURN STD_LOGIC_VECTOR;
---
FUNCTION LIMPIAR_PANTALLA(DATO9 : STD_LOGIC)RETURN STD_LOGIC_VECTOR;

CONSTANT a:INTEGER:=1;CONSTANT j:INTEGER:=10;CONSTANT s:INTEGER:=19;
CONSTANT b:INTEGER:=2;CONSTANT k:INTEGER:=11;CONSTANT t:INTEGER:=20;
CONSTANT c:INTEGER:=3;CONSTANT l:INTEGER:=12;CONSTANT u:INTEGER:=21;
CONSTANT d:INTEGER:=4;CONSTANT m:INTEGER:=13;CONSTANT v:INTEGER:=22;
CONSTANT e:INTEGER:=5;CONSTANT n:INTEGER:=14;CONSTANT w:INTEGER:=23;
CONSTANT f:INTEGER:=6;CONSTANT o:INTEGER:=15;CONSTANT x:INTEGER:=24;
CONSTANT g:INTEGER:=7;CONSTANT p:INTEGER:=16;CONSTANT y:INTEGER:=25;
CONSTANT h:INTEGER:=8;CONSTANT q:INTEGER:=17;CONSTANT z:INTEGER:=26;
CONSTANT i:INTEGER:=9;CONSTANT r:INTEGER:=18;

CONSTANT Ma:INTEGER:=27;CONSTANT Mj:INTEGER:=36;CONSTANT MAs:INTEGER:=45;
CONSTANT Mb:INTEGER:=28;CONSTANT Mk:INTEGER:=37;CONSTANT Mt:INTEGER:=46;
CONSTANT Mc:INTEGER:=29;CONSTANT Ml:INTEGER:=38;CONSTANT Mu:INTEGER:=47;
CONSTANT Md:INTEGER:=30;CONSTANT Mm:INTEGER:=39;CONSTANT Mv:INTEGER:=48;
CONSTANT Me:INTEGER:=31;CONSTANT Mn:INTEGER:=40;CONSTANT Mw:INTEGER:=49;
CONSTANT Mf:INTEGER:=32;CONSTANT Mo:INTEGER:=41;CONSTANT Mx:INTEGER:=50;
CONSTANT Mg:INTEGER:=33;CONSTANT Mp:INTEGER:=42;CONSTANT My:INTEGER:=51;
CONSTANT Mh:INTEGER:=34;CONSTANT Mq:INTEGER:=43;CONSTANT Mz:INTEGER:=52;
CONSTANT Mi:INTEGER:=35;CONSTANT Mr:INTEGER:=44;

end COMANDOS_LCDSPI_REVA;


package body COMANDOS_LCDSPI_REVA is

----LCD_INI()------
-------------------
FUNCTION LCD_INI(DATO : STD_LOGIC_VECTOR(1 DOWNTO 0)) RETURN STD_LOGIC_VECTOR IS
VARIABLE DATAOUT : STD_LOGIC_VECTOR(11 DOWNTO 0);
BEGIN
CASE DATO IS
WHEN "00" => RETURN x"101";
WHEN "01" => RETURN x"102";
WHEN "10" => RETURN x"103";
WHEN OTHERS => RETURN x"104";
END CASE;
END LCD_INI;
-----------------

-----CHAR()-----
-----------------
FUNCTION CHAR(DATO1 : INTEGER) RETURN STD_LOGIC_VECTOR IS
VARIABLE DATAOUT1 : STD_LOGIC_VECTOR(11 DOWNTO 0);
BEGIN
CASE DATO1 IS
WHEN 1 => RETURN x"109";
WHEN 2 => RETURN x"10A";
WHEN 3 => RETURN x"10B";
WHEN 4 => RETURN x"10C";
WHEN 5 => RETURN x"10D";
WHEN 6 => RETURN x"10E";
WHEN 7 => RETURN x"10F";
WHEN 8 => RETURN x"110";
WHEN 9 => RETURN x"111";
WHEN 10 => RETURN x"112";
WHEN 11 => RETURN x"113";
WHEN 12 => RETURN x"114";
WHEN 13 => RETURN x"115";
WHEN 14 => RETURN x"116";
WHEN 15 => RETURN x"117";
WHEN 16 => RETURN x"118";
WHEN 17 => RETURN x"119";
WHEN 18 => RETURN x"11A";
WHEN 19 => RETURN x"11B";
WHEN 20 => RETURN x"11C";
WHEN 21 => RETURN x"11D";
WHEN 22 => RETURN x"11E";
WHEN 23 => RETURN x"11F";
WHEN 24 => RETURN x"120";
WHEN 25 => RETURN x"121";
WHEN 26 => RETURN x"122";
----
WHEN 27 => RETURN x"123";
WHEN 28 => RETURN x"124";
WHEN 29 => RETURN x"125";
WHEN 30 => RETURN x"126";
WHEN 31 => RETURN x"127";
WHEN 32 => RETURN x"128";
WHEN 33 => RETURN x"129";
WHEN 34 => RETURN x"12A";
WHEN 35 => RETURN x"12B";
WHEN 36 => RETURN x"12C";
WHEN 37 => RETURN x"12D";
WHEN 38 => RETURN x"12E";
WHEN 39 => RETURN x"12F";
WHEN 40 => RETURN x"130";
WHEN 41 => RETURN x"131";
WHEN 42 => RETURN x"132";
WHEN 43 => RETURN x"133";
WHEN 44 => RETURN x"134";
WHEN 45 => RETURN x"135";
WHEN 46 => RETURN x"136";
WHEN 47 => RETURN x"137";
WHEN 48 => RETURN x"138";
WHEN 49 => RETURN x"139";
WHEN 50 => RETURN x"13A";
WHEN 51 => RETURN x"13B";
WHEN 52 => RETURN x"13C";
----
WHEN OTHERS => RETURN x"147";
END CASE;
END CHAR;
  
---INT_NUM()----
----------------

FUNCTION INT_NUM(DATO10 : INTEGER) RETURN STD_LOGIC_VECTOR IS
VARIABLE DATAOUT6 : STD_LOGIC_VECTOR(11 DOWNTO 0);
BEGIN
CASE DATO10 IS
WHEN 0 => RETURN x"030";
WHEN 1 => RETURN x"031";
WHEN 2 => RETURN x"032";
WHEN 3 => RETURN x"033";
WHEN 4 => RETURN x"034";
WHEN 5 => RETURN x"035";
WHEN 6 => RETURN x"036";
WHEN 7 => RETURN x"037";
WHEN 8 => RETURN x"038";
WHEN 9 => RETURN x"039";
WHEN OTHERS => RETURN x"030";
END CASE;
END INT_NUM;

----------------
  
----POS()------
--------------------
FUNCTION POS(DATO2,DATO3 : INTEGER) RETURN STD_LOGIC_VECTOR IS
VARIABLE DATAOUT2 : STD_LOGIC_VECTOR(11 DOWNTO 0);
BEGIN
IF 	DATO2 = 1 AND DATO3 = 1  THEN RETURN x"150";
ELSIF DATO2 = 1 AND DATO3 = 2  THEN RETURN x"151";
ELSIF DATO2 = 1 AND DATO3 = 3  THEN RETURN x"152";
ELSIF DATO2 = 1 AND DATO3 = 4  THEN RETURN x"153";
ELSIF DATO2 = 1 AND DATO3 = 5  THEN RETURN x"154";
ELSIF DATO2 = 1 AND DATO3 = 6  THEN RETURN x"155";
ELSIF DATO2 = 1 AND DATO3 = 7  THEN RETURN x"156";
ELSIF DATO2 = 1 AND DATO3 = 8  THEN RETURN x"157";
ELSIF DATO2 = 1 AND DATO3 = 9  THEN RETURN x"158";
ELSIF DATO2 = 1 AND DATO3 = 10 THEN RETURN x"159";
ELSIF DATO2 = 1 AND DATO3 = 11 THEN RETURN x"15A";
ELSIF DATO2 = 1 AND DATO3 = 12 THEN RETURN x"15B";
ELSIF DATO2 = 1 AND DATO3 = 13 THEN RETURN x"15C";
ELSIF DATO2 = 1 AND DATO3 = 14 THEN RETURN x"15D";
ELSIF DATO2 = 1 AND DATO3 = 15 THEN RETURN x"15E";
ELSIF DATO2 = 1 AND DATO3 = 16 THEN RETURN x"15F";
ELSIF DATO2 = 1 AND DATO3 = 17 THEN RETURN x"160";
ELSIF DATO2 = 1 AND DATO3 = 18 THEN RETURN x"161";
ELSIF DATO2 = 1 AND DATO3 = 19 THEN RETURN x"162";
ELSIF DATO2 = 1 AND DATO3 = 20 THEN RETURN x"163";
-------
ELSIF	DATO2 = 2 AND DATO3 = 1  THEN RETURN x"164";
ELSIF DATO2 = 2 AND DATO3 = 2  THEN RETURN x"165";
ELSIF DATO2 = 2 AND DATO3 = 3  THEN RETURN x"166";
ELSIF DATO2 = 2 AND DATO3 = 4  THEN RETURN x"167";
ELSIF DATO2 = 2 AND DATO3 = 5  THEN RETURN x"168";
ELSIF DATO2 = 2 AND DATO3 = 6  THEN RETURN x"169";
ELSIF DATO2 = 2 AND DATO3 = 7  THEN RETURN x"16A";
ELSIF DATO2 = 2 AND DATO3 = 8  THEN RETURN x"16B";
ELSIF DATO2 = 2 AND DATO3 = 9  THEN RETURN x"16C";
ELSIF DATO2 = 2 AND DATO3 = 10 THEN RETURN x"16D";
ELSIF DATO2 = 2 AND DATO3 = 11 THEN RETURN x"16E";
ELSIF DATO2 = 2 AND DATO3 = 12 THEN RETURN x"16F";
ELSIF DATO2 = 2 AND DATO3 = 13 THEN RETURN x"170";
ELSIF DATO2 = 2 AND DATO3 = 14 THEN RETURN x"171";
ELSIF DATO2 = 2 AND DATO3 = 15 THEN RETURN x"172";
ELSIF DATO2 = 2 AND DATO3 = 16 THEN RETURN x"173";
ELSIF DATO2 = 2 AND DATO3 = 17 THEN RETURN x"174";
ELSIF DATO2 = 2 AND DATO3 = 18 THEN RETURN x"175";
ELSIF DATO2 = 2 AND DATO3 = 19 THEN RETURN x"176";
ELSIF DATO2 = 2 AND DATO3 = 20 THEN RETURN x"177";
ELSE RETURN x"177";
--ELSE NULL;
END IF;
END POS;
-------------------

------BUCLE_INI()----
----------------------
FUNCTION BUCLE_INI(DATO8 : INTEGER)RETURN STD_LOGIC_VECTOR IS
VARIABLE DATAOUT6 : STD_LOGIC_VECTOR(11 DOWNTO 0);
BEGIN
IF DATO8 = 1 THEN RETURN x"17C";
ELSE RETURN x"17C";
END IF;
END BUCLE_INI;
-------------------

------BUCLE_FIN()----
----------------------
FUNCTION BUCLE_FIN(DATO9 : INTEGER)RETURN STD_LOGIC_VECTOR IS
VARIABLE DATAOUT7 : STD_LOGIC_VECTOR(11 DOWNTO 0);
BEGIN
IF DATO9 = 1 THEN RETURN x"17D";
ELSE RETURN x"17D";
END IF;
END BUCLE_FIN;
-------------------

------LIMPIAR_PANTALLA()----
----------------------
FUNCTION LIMPIAR_PANTALLA(DATO9 : STD_LOGIC)RETURN STD_LOGIC_VECTOR IS
VARIABLE DATAOUT10 : STD_LOGIC_VECTOR(11 DOWNTO 0);
BEGIN
IF DATO9 = '1' THEN RETURN x"1FE";
ELSE RETURN x"1FD";
END IF;
END LIMPIAR_PANTALLA;
-------------------


------CHAR_ASCII()----
----------------------
FUNCTION CHAR_ASCII(DATO6 : STD_LOGIC_VECTOR(7 DOWNTO 0))RETURN STD_LOGIC_VECTOR IS
VARIABLE DATAOUT4 : STD_LOGIC_VECTOR(11 DOWNTO 0);
BEGIN
DATAOUT4 := "0000"&DATO6;
RETURN DATAOUT4;

END CHAR_ASCII;
-------------------


------CODIGO_FIN()----
----------------------
FUNCTION CODIGO_FIN(DATO7 : INTEGER)RETURN STD_LOGIC_VECTOR IS
VARIABLE DATAOUT5 : STD_LOGIC_VECTOR(11 DOWNTO 0);
BEGIN
IF DATO7 = 1 THEN RETURN x"1FF";
ELSE RETURN x"1FF";
END IF;
END CODIGO_FIN;
-------------------

 
end COMANDOS_LCDSPI_REVA;
